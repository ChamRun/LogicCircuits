// Verilog Test Fixture Template

  `timescale 1 ns / 1 ps

  module TEST_gate;
          
   initial begin
      $display("\n\nMy String\n\n");
   end

  endmodule
