`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:57:20 11/17/2021 
// Design Name: 
// Module Name:    mux_four_one 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module mux_tb();

	 wire out;
    reg w3, w2, w1, w0, s1, s0;
     
    always begin
	
		#1 w3 = 0; w2 = 0; w1 = 0; w0 = 0; s1 = 0; s0 = 0;
		#1 w3 = 0; w2 = 0; w1 = 0; w0 = 0; s1 = 0; s0 = 1;
		#1 w3 = 0; w2 = 0; w1 = 0; w0 = 0; s1 = 1; s0 = 0;
		#1 w3 = 0; w2 = 0; w1 = 0; w0 = 0; s1 = 1; s0 = 1;
		
		#1 w3 = 0; w2 = 0; w1 = 0; w0 = 1; s1 = 0; s0 = 0;
		#1 w3 = 0; w2 = 0; w1 = 0; w0 = 1; s1 = 0; s0 = 1;
		#1 w3 = 0; w2 = 0; w1 = 0; w0 = 1; s1 = 1; s0 = 0;
		#1 w3 = 0; w2 = 0; w1 = 0; w0 = 1; s1 = 1; s0 = 1;
		
		#1 w3 = 0; w2 = 0; w1 = 1; w0 = 0; s1 = 0; s0 = 0;
		#1 w3 = 0; w2 = 0; w1 = 1; w0 = 0; s1 = 0; s0 = 1;
		#1 w3 = 0; w2 = 0; w1 = 1; w0 = 0; s1 = 1; s0 = 0;
		#1 w3 = 0; w2 = 0; w1 = 1; w0 = 0; s1 = 1; s0 = 1;
		
		#1 w3 = 0; w2 = 0; w1 = 1; w0 = 1; s1 = 0; s0 = 0;
		#1 w3 = 0; w2 = 0; w1 = 1; w0 = 1; s1 = 0; s0 = 1;
		#1 w3 = 0; w2 = 0; w1 = 1; w0 = 1; s1 = 1; s0 = 0;
		#1 w3 = 0; w2 = 0; w1 = 1; w0 = 1; s1 = 1; s0 = 1;
		
		#1 w3 = 0; w2 = 1; w1 = 0; w0 = 0; s1 = 0; s0 = 0;
		#1 w3 = 0; w2 = 1; w1 = 0; w0 = 0; s1 = 0; s0 = 1;
		#1 w3 = 0; w2 = 1; w1 = 0; w0 = 0; s1 = 1; s0 = 0;
		#1 w3 = 0; w2 = 1; w1 = 0; w0 = 0; s1 = 1; s0 = 1;
		
		#1 w3 = 0; w2 = 1; w1 = 0; w0 = 1; s1 = 0; s0 = 0;
		#1 w3 = 0; w2 = 1; w1 = 0; w0 = 1; s1 = 0; s0 = 1;
		#1 w3 = 0; w2 = 1; w1 = 0; w0 = 1; s1 = 1; s0 = 0;
		#1 w3 = 0; w2 = 1; w1 = 0; w0 = 1; s1 = 1; s0 = 1;
		
		#1 w3 = 0; w2 = 1; w1 = 1; w0 = 0; s1 = 0; s0 = 0;
		#1 w3 = 0; w2 = 1; w1 = 1; w0 = 0; s1 = 0; s0 = 1;
		#1 w3 = 0; w2 = 1; w1 = 1; w0 = 0; s1 = 1; s0 = 0;
		#1 w3 = 0; w2 = 1; w1 = 1; w0 = 0; s1 = 1; s0 = 1;
		
		#1 w3 = 0; w2 = 1; w1 = 1; w0 = 1; s1 = 0; s0 = 0;
		#1 w3 = 0; w2 = 1; w1 = 1; w0 = 1; s1 = 0; s0 = 1;
		#1 w3 = 0; w2 = 1; w1 = 1; w0 = 1; s1 = 1; s0 = 0;
		#1 w3 = 0; w2 = 1; w1 = 1; w0 = 1; s1 = 1; s0 = 1;
		
		
		
		#1 w3 = 1; w2 = 0; w1 = 0; w0 = 0; s1 = 0; s0 = 0;
		#1 w3 = 1; w2 = 0; w1 = 0; w0 = 0; s1 = 0; s0 = 1;
		#1 w3 = 1; w2 = 0; w1 = 0; w0 = 0; s1 = 1; s0 = 0;
		#1 w3 = 1; w2 = 0; w1 = 0; w0 = 0; s1 = 1; s0 = 1;
		
		#1 w3 = 1; w2 = 0; w1 = 0; w0 = 1; s1 = 0; s0 = 0;
		#1 w3 = 1; w2 = 0; w1 = 0; w0 = 1; s1 = 0; s0 = 1;
		#1 w3 = 1; w2 = 0; w1 = 0; w0 = 1; s1 = 1; s0 = 0;
		#1 w3 = 1; w2 = 0; w1 = 0; w0 = 1; s1 = 1; s0 = 1;
		
		#1 w3 = 1; w2 = 0; w1 = 1; w0 = 0; s1 = 0; s0 = 0;
		#1 w3 = 1; w2 = 0; w1 = 1; w0 = 0; s1 = 0; s0 = 1;
		#1 w3 = 1; w2 = 0; w1 = 1; w0 = 0; s1 = 1; s0 = 0;
		#1 w3 = 1; w2 = 0; w1 = 1; w0 = 0; s1 = 1; s0 = 1;
		
		#1 w3 = 1; w2 = 0; w1 = 1; w0 = 1; s1 = 0; s0 = 0;
		#1 w3 = 1; w2 = 0; w1 = 1; w0 = 1; s1 = 0; s0 = 1;
		#1 w3 = 1; w2 = 0; w1 = 1; w0 = 1; s1 = 1; s0 = 0;
		#1 w3 = 1; w2 = 0; w1 = 1; w0 = 1; s1 = 1; s0 = 1;
	
		#1 w3 = 1; w2 = 1; w1 = 0; w0 = 0; s1 = 0; s0 = 0;
		#1 w3 = 1; w2 = 1; w1 = 0; w0 = 0; s1 = 0; s0 = 1;
		#1 w3 = 1; w2 = 1; w1 = 0; w0 = 0; s1 = 1; s0 = 0;
		#1 w3 = 1; w2 = 1; w1 = 0; w0 = 0; s1 = 1; s0 = 1;
		
		#1 w3 = 1; w2 = 1; w1 = 0; w0 = 1; s1 = 0; s0 = 0;
		#1 w3 = 1; w2 = 1; w1 = 0; w0 = 1; s1 = 0; s0 = 1;
		#1 w3 = 1; w2 = 1; w1 = 0; w0 = 1; s1 = 1; s0 = 0;
		#1 w3 = 1; w2 = 1; w1 = 0; w0 = 1; s1 = 1; s0 = 1;
		
		#1 w3 = 1; w2 = 1; w1 = 1; w0 = 0; s1 = 0; s0 = 0;
		#1 w3 = 1; w2 = 1; w1 = 1; w0 = 0; s1 = 0; s0 = 1;
		#1 w3 = 1; w2 = 1; w1 = 1; w0 = 0; s1 = 1; s0 = 0;
		#1 w3 = 1; w2 = 1; w1 = 1; w0 = 0; s1 = 1; s0 = 1;
		
		#1 w3 = 1; w2 = 1; w1 = 1; w0 = 1; s1 = 0; s0 = 0;
		#1 w3 = 1; w2 = 1; w1 = 1; w0 = 1; s1 = 0; s0 = 1;
		#1 w3 = 1; w2 = 1; w1 = 1; w0 = 1; s1 = 1; s0 = 0;
		#1 w3 = 1; w2 = 1; w1 = 1; w0 = 1; s1 = 1; s0 = 1;
	 
	 end
     
    initial begin
		//Initialize clock
		w3 = 0;
		w2 = 0;
		w1 = 0;
		w0 = 0;
		s1 = 0;
		s0 = 0;
     
		//End simulation
		#65
		$finish;
    end
     
	 mux_four_one myGate(out, w3, w2, w1, w0, s1, s0);
	 
endmodule



module mux_four_one(y, w3, w2, w1, w0, s1, s0);

	input w0, w1, w2, w3;
	input s0, s1;
	output y;
	
	wire not_s0, not_s1;
	not g0(not_s0, s0),
		 g1(not_s1, s1);
		 
	
	wire a, b, c, d;
	and g2(a, w0, not_s1, not_s0),
		 g3(b, w1, not_s1, s0),
		 g4(c, w2, s1, not_s0),
		 g5(d, w3, s1, s0);
		 
	or g6(y, a, b, c, d);
	

endmodule

